LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY divf IS
	GENERIC(FREC: INTEGER := 24999); -- FREC = (50 MHz/2*Fdeseada) - 1
	-- 24999    >> 1 kHz
	-- 249999   >> 100 Hz
	-- 24999999 >> 1 Hz
	PORT(CLK_MST: IN STD_LOGIC; -- RELOJ PRINCIPAL
			   CLK: BUFFER STD_LOGIC);
END ENTITY;

ARCHITECTURE BEAS OF divf IS
SIGNAL AUX: INTEGER RANGE 0 TO FREC;
BEGIN
	PROCESS(CLK_MST)
	BEGIN
		IF RISING_EDGE (CLK_MST) THEN
			IF AUX = 0 THEN
				CLK <= NOT CLK;
				AUX <= FREC;
			ELSE
				AUX <= AUX - 1;
			END IF;
		END IF;
	END PROCESS;

END BEAS;