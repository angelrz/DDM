LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ram IS
PORT(CLK, RW:STD_LOGIC;
			DIR: IN INTEGER RANGE 0 TO 3;
			DATO: IN INTEGER RANGE 0 TO 15;
			SAL: OUT INTEGER RANGE 0 TO 15);

END ENTITY;
ARCHITECTURE BEAS OF ram IS
TYPE MEMORIA IS ARRAY (0 TO 3) OF INTEGER RANGE 0 TO 15; -- ARREGLO DE N DE 8 BITS.
SIGNAL ADDR: MEMORIA;
	BEGIN
	PROCESS(CLK)
	BEGIN
		IF RISING_EDGE (CLK) THEN
			IF RW='1' THEN -- ESCRIBRIR
				ADDR(DIR) <= DATO;
			ELSE -- LEER
				SAL <= ADDR(DIR);
			END IF;
		END IF;
	END PROCESS;
END BEAS;