LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY deco_num IS
PORT(NUM: in INTEGER RANGE 0 to 7;
		SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END deco_num;

ARCHITECTURE am OF deco_num IS
	BEGIN
	WITH NUM SELECT
	-- Decodificador de 1-7
	SEG <= "00000011" WHEN 0,
			 "10011111" WHEN 1,
			 "00100101" WHEN 2,
			 "00001101" WHEN 3,
			 "10011001" WHEN 4,
			 "01001001" WHEN 5,
			 "01000001" WHEN 6,
			 "00011101" WHEN OTHERS;
end am;