LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY deco_let IS
	PORT(NUM: in INTEGER RANGE 0 to 7;
		SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END deco_let;

ARCHITECTURE am OF deco_let IS
	BEGIN
	WITH NUM SELECT
	SEG <= "00010001" WHEN 0,
			 "11000001" WHEN 1,
			 "01100011" WHEN 2,
			 "10000101" WHEN 3,
			 "01100001" WHEN 4,
			 "01110001" WHEN 5,
			 "00001001" WHEN 6,
			 "10010001" WHEN 7;
END am;